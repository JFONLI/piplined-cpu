module Imm_Gen(
    data_i,
    data_o
    );

//I/O ports
input   [32-1:0] data_i;
output  [64-1:0] data_o;

//Internal Signals
reg     [64-1:0] data_o;

//Gen Imm

endmodule